library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--------------------------------------------------
package componentsRISC is
	
	component dregister is --tested
	port (DIN: in std_logic_vector(15 downto 0); 
		  clk, en: in std_logic; 
		  DOUT: out std_logic_vector(15 downto 0));
	end component;
	
	component dflipflop is --tested
	port (DIN: in std_logic; 
		  clk, en: in std_logic; 
		  DOUT: out std_logic);
	end component;
	
	component mux2_16 is --tested
	port (IN1,IN0: in std_logic_vector(15 downto 0); 
		  s: in std_logic; 
		  OUTPUT: out std_logic_vector(15 downto 0));
	end component;
	
	component mux4_16 is --tested
	port (IN3,IN2,IN1,IN0: in std_logic_vector(15 downto 0); 
		  s: in std_logic_vector(1 downto 0); 
		  OUTPUT: out std_logic_vector(15 downto 0));
	end component;
	
	component mux8_16 is --tested
	port (IN7,IN6,IN5,IN4,IN3,IN2,IN1,IN0: in std_logic_vector(15 downto 0); 
		  s: in std_logic_vector(2 downto 0); 
		  OUTPUT: out std_logic_vector(15 downto 0));
	end component;
	
	component mux2_3 is --tested
	port (IN1,IN0: in std_logic_vector(2 downto 0); 
		  s: in std_logic; 
		  OUTPUT: out std_logic_vector(2 downto 0));
	end component;
	
	component mux4_3 is --tested
	port (IN3,IN2,IN1,IN0: in std_logic_vector(2 downto 0); 
		  s: in std_logic_vector(1 downto 0); 
		  OUTPUT: out std_logic_vector(2 downto 0));
	end component;
	
	component mux8_3 is --tested
	port (IN7,IN6,IN5,IN4,IN3,IN2,IN1,IN0: in std_logic_vector(2 downto 0); 
		  s: in std_logic_vector(2 downto 0); 
		  OUTPUT: out std_logic_vector(2 downto 0));
	end component;
	
	component priority is --tested
	port (INPUT: in std_logic_vector(8 downto 0); 
		  output: out std_logic_vector(2 downto 0); 
		  valid: out std_logic);
	end component;

	component ir_decoder is
	port (s: in std_logic_vector(2 downto 0); 
		  IR: in std_logic_vector(15 downto 0); 
		  new_IR: out std_logic_vector(15 downto 0));
	end component;

	component register_file is
	port (
		   a1,a2,a3: in std_logic_vector(2 downto 0);   --a3 is the address where data to be written , a2 a1 to read the data
		   d3: in std_logic_vector(15 downto 0);        -- d3 is the daata to write 
			wr: in std_logic;                            
			d1, d2: out std_logic_vector(15 downto 0);
			reset: in std_logic;
			clk: in std_logic);
	end component;
	
	component LeftShift is 
	port (IN1: in std_logic_vector(8 downto 0); 
		  OUTPUT1: out std_logic_vector(15 downto 0));
	end component;
	
	component SgnExtd7 is 
	port (IN1: in std_logic_vector(8 downto 0); 
		  OUTPUT1: out std_logic_vector(15 downto 0));
	end component;
	
	component SgnExtd10 is 
	port (IN1: in std_logic_vector(5 downto 0); 
		  OUTPUT1: out std_logic_vector(15 downto 0));
	end component;

	component memory is --tested
    generic (data_width: integer:= 16; addr_width: integer := 16);
    port(din: in std_logic_vector(data_width-1 downto 0);
        dout: out std_logic_vector(data_width-1 downto 0);
        rbar: in std_logic;
        wbar: in std_logic;
        addrin: in std_logic_vector(addr_width-1 downto 0));
	end component;
	
	component alu is 
	port( X,Y : in std_logic_vector(15 downto 0); 
		  op_code_bits : in std_logic_vector(3 downto 0); 
		  cz_bits : in std_logic_vector(1 downto 0);
		  OUTPUT_ALU : out std_logic_vector(15 downto 0);
		  carry_ALU,zero_ALU : out std_logic);
	end component;
	
end package;
---------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity dregister is                  -- no. of bits
  port (
    din  : in  std_logic_vector(15 downto 0);
    dout : out std_logic_vector(15 downto 0);
    en: in std_logic;
    clk     : in  std_logic);
end dregister;

architecture behave of dregister is

begin  -- behave
process(clk)
begin 
  if(clk'event and clk = '1') then
    if en = '1' then
      dout <= din;
    end if;
  end if;
end process;
end behave;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity dflipflop is                  -- no. of bits
  port (
    din  : in  std_logic;
    dout : out std_logic;
    en: in std_logic;
    clk     : in std_logic);
end dflipflop;

architecture behave of dflipflop is

begin  -- behave
process(clk)
begin 
  if(clk'event and clk = '1') then
    if en = '1' then
      dout <= din;
    end if;
  end if;
end process;
end behave;
-----------------------------------------------------------
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity mux2_16 is
	port (IN1,IN0: in std_logic_vector(15 downto 0); s: in std_logic; OUTPUT: out std_logic_vector(15 downto 0));
end mux2_16;

architecture behave_mux2_16 of mux2_16 is
begin
process(s, IN0, IN1)
begin
	if(s='0') then OUTPUT <= IN0;
	end if;
	if(s='1') then OUTPUT <= IN1;
	end if;
end process;
end behave_mux2_16;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity mux4_16 is
	port (IN3,IN2,IN1,IN0: in std_logic_vector(15 downto 0); s: in std_logic_vector(1 downto 0); OUTPUT: out std_logic_vector(15 downto 0));
end mux4_16;

architecture behave_mux4_16 of mux4_16 is
begin
process(s, IN0, IN1, IN2, IN3)
begin
	if(s="00") then OUTPUT <= IN0;
	end if;
	if(s="01") then OUTPUT <= IN1;
	end if;
	if(s="10") then OUTPUT <= IN2;
	end if;
	if(s="11") then OUTPUT <= IN3;
	end if;
end process;
end behave_mux4_16;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity mux8_16 is
	port (IN7,IN6,IN5,IN4,IN3,IN2,IN1,IN0: in std_logic_vector(15 downto 0); s: in std_logic_vector(2 downto 0); OUTPUT: out std_logic_vector(15 downto 0));
end mux8_16;

architecture behave_mux8_16 of mux8_16 is
begin
process(s, IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7)
begin
	if(s="000") then OUTPUT <= IN0;
	end if;
	if(s="001") then OUTPUT <= IN1;
	end if;
	if(s="010") then OUTPUT <= IN2;
	end if;
	if(s="011") then OUTPUT <= IN3;
	end if;
	if(s="100") then OUTPUT <= IN4;
	end if;
	if(s="101") then OUTPUT <= IN5;
	end if;
	if(s="110") then OUTPUT <= IN6;
	end if;
	if(s="111") then OUTPUT <= IN7;
	end if;
end process;
end behave_mux8_16;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;


entity mux2_3 is
	port (IN1,IN0: in std_logic_vector(2 downto 0); s: in std_logic; OUTPUT: out std_logic_vector(2 downto 0));
end mux2_3;

architecture behave_mux2_3 of mux2_3 is
begin
process(s, IN0, IN1)
begin
	if(s='0') then OUTPUT <= IN0;
	end if;
	if(s='1') then OUTPUT <= IN1;
	end if;
end process;
end behave_mux2_3;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity mux4_3 is
	port (IN3,IN2,IN1,IN0: in std_logic_vector(2 downto 0); s: in std_logic_vector(1 downto 0); OUTPUT: out std_logic_vector(2 downto 0));
end mux4_3;

architecture behave_mux4_3 of mux4_3 is
begin
process(s, IN0, IN1, IN2, IN3)
begin
	if(s="00") then OUTPUT <= IN0;
	end if;
	if(s="01") then OUTPUT <= IN1;
	end if;
	if(s="10") then OUTPUT <= IN2;
	end if;
	if(s="11") then OUTPUT <= IN3;
	end if;
end process;
end behave_mux4_3;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity mux8_3 is
	port (IN7,IN6,IN5,IN4,IN3,IN2,IN1,IN0: in std_logic_vector(2 downto 0); s: in std_logic_vector(2 downto 0); OUTPUT: out std_logic_vector(2 downto 0));
end mux8_3;

architecture behave_mux8_3 of mux8_3 is
begin
process(s, IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7)
begin
	if(s="000") then OUTPUT <= IN0;
	end if;
	if(s="001") then OUTPUT <= IN1;
	end if;
	if(s="010") then OUTPUT <= IN2;
	end if;
	if(s="011") then OUTPUT <= IN3;
	end if;
	if(s="100") then OUTPUT <= IN4;
	end if;
	if(s="101") then OUTPUT <= IN5;
	end if;
	if(s="110") then OUTPUT <= IN6;
	end if;
	if(s="111") then OUTPUT <= IN7;
	end if;
end process;
end behave_mux8_3;
-----------------------------------------------------------








library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity priority is
	port (INPUT: in std_logic_vector(8 downto 0); output: out std_logic_vector(2 downto 0); valid: out std_logic);
	end priority; 

architecture behave_priority of priority is
begin
process(INPUT)
begin
	if (INPUT(0)='1') then OUTPUT <= "000";
	elsif (INPUT(1)='1') then OUTPUT <= "001";
	elsif (INPUT(2)='1') then OUTPUT <= "010";
	elsif (INPUT(3)='1') then OUTPUT <= "011";
	elsif (INPUT(4)='1') then OUTPUT <= "100";
	elsif (INPUT(5)='1') then OUTPUT <= "101";
	elsif (INPUT(6)='1') then OUTPUT <= "110";
	elsif (INPUT(7)='1') then OUTPUT <= "111";
	else OUTPUT <= "000";
	end if;
	if (INPUT="000000000") then valid <= '0';
	else valid <= '1';
	end if;
end process;
end behave_priority;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity ir_decoder is
	port (s: in std_logic_vector(2 downto 0); IR: in std_logic_vector(15 downto 0); new_IR: out std_logic_vector(15 downto 0));
end ir_decoder;

architecture behave_ir_dec of ir_decoder is
signal temp: std_logic_vector(15 downto 0);
begin
process(s, IR, temp)
begin
	if(s="000") then temp(0) <= '1'; end if;
	if(s="001") then temp(1) <= '1'; end if;
	if(s="010") then temp(2) <= '1'; end if;
	if(s="011") then temp(3) <= '1'; end if;
	if(s="100") then temp(4) <= '1'; end if;
	if(s="101") then temp(5) <= '1'; end if;
	if(s="110") then temp(6) <= '1'; end if;
	if(s="111") then temp(7) <= '1'; end if;
	temp(15 downto 8) <= "00000000";
	new_IR <= IR xor temp;
end process;
end behave_ir_dec;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_bit.all;

entity register_file is
	port (
	a1,a2,a3: in std_logic_vector(2 downto 0);   --a3 is the address where data to be written , a2 a1 to read the data
	d3: in std_logic_vector(15 downto 0);        -- d3 is the daata to write 
	wr: in std_logic;                            
	d1, d2: out std_logic_vector(15 downto 0);
	reset: in std_logic;
	clk: in std_logic
	);
end entity register_file;

architecture behave_rf of register_file is
  type registerFile is array(0 to 7) of std_logic_vector(15 downto 0);
  signal registers : registerFile;
  
  function To_Integer(x: bit_vector) return integer is
      variable xu: unsigned(x'range);
   begin
      for I in x'range loop
         xu(I) := x(I);
      end loop;
      return(To_Integer(xu));
   end To_Integer;

   function to_bit_vector(x: std_logic_vector) return bit_vector is
      variable ret_val: bit_vector(1 to x'length);
      alias lx: std_logic_vector(1 to x'length) is x;
  begin
 	for I in 1 to x'length loop
		if(lx(I) = '1') then
			ret_val(I) := '1';
		else
			ret_val(I) := '0';
		end if;
	end loop;
	return(ret_val);
  end to_bit_vector;
  
begin
  regFile : process (clk,wr,a1,a2,a3,d3,reset) is
  begin      
	if (reset='1') then
		registers(7) <= "0000000000000000";
	else
		if (clk'event and clk = '1') then
			if wr='1' then
				registers(to_Integer(to_bit_vector(a3))) <= d3;  -- Write
			end if;
		end if;
		d1 <= registers(to_Integer(to_bit_vector(a1)));
		d2 <= registers(to_Integer(to_bit_vector(a2))); 
	end if;
  end process;
end behave_rf;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity LeftShift is 
	port (IN1: in std_logic_vector(8 downto 0); OUTPUT1: out std_logic_vector(15 downto 0));
end LeftShift;

architecture behave_LeftShift of LeftShift is
begin
process(IN1)
begin
	OUTPUT1(0) <= '0';
	OUTPUT1(1) <= '0';
	OUTPUT1(2) <= '0';
	OUTPUT1(3) <= '0';
	OUTPUT1(4) <= '0';
	OUTPUT1(5) <= '0';
	OUTPUT1(6) <= '0';
	OUTPUT1(7) <= IN1(0);
	OUTPUT1(8) <= IN1(1);
	OUTPUT1(9) <= IN1(2);
	OUTPUT1(10) <= IN1(3);
	OUTPUT1(11) <= IN1(4);
	OUTPUT1(12) <= IN1(5);
	OUTPUT1(13) <= IN1(6);
	OUTPUT1(14) <= IN1(7);
	OUTPUT1(15) <= IN1(8);
end process;
end behave_LeftShift;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity SgnExtd7 is 
	port (IN1: in std_logic_vector(8 downto 0); OUTPUT1: out std_logic_vector(15 downto 0));
end SgnExtd7;

architecture behave_SgnExtd7 of SgnExtd7 is
begin
process(IN1)
begin
	OUTPUT1(0) <= IN1(0);
	OUTPUT1(1) <= IN1(1);
	OUTPUT1(2) <= IN1(2);
	OUTPUT1(3) <= IN1(3);
	OUTPUT1(4) <= IN1(4);
	OUTPUT1(5) <= IN1(5);
	OUTPUT1(6) <= IN1(6);
	OUTPUT1(7) <= IN1(7);
	OUTPUT1(8) <= IN1(8);
	OUTPUT1(9) <= IN1(8);
	OUTPUT1(10) <= IN1(8);
	OUTPUT1(11) <= IN1(8);
	OUTPUT1(12) <= IN1(8);
	OUTPUT1(13) <= IN1(8);
	OUTPUT1(14) <= IN1(8);
	OUTPUT1(15) <= IN1(8);

end process;
end behave_SgnExtd7;
-----------------------------------------------------------

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

entity SgnExtd10 is 
	port (IN1: in std_logic_vector(5 downto 0); OUTPUT1: out std_logic_vector(15 downto 0));
end SgnExtd10;

architecture behave_SgnExtd10 of SgnExtd10 is
begin
process(IN1)
begin
	OUTPUT1(0) <= IN1(0);
	OUTPUT1(1) <= IN1(1);
	OUTPUT1(2) <= IN1(2);
	OUTPUT1(3) <= IN1(3);
	OUTPUT1(4) <= IN1(4);
	OUTPUT1(5) <= IN1(5);
	OUTPUT1(6) <= IN1(5);
	OUTPUT1(7) <= IN1(5);
	OUTPUT1(8) <= IN1(5);
	OUTPUT1(9) <= IN1(5);
	OUTPUT1(10) <= IN1(5);
	OUTPUT1(11) <= IN1(5);
	OUTPUT1(12) <= IN1(5);
	OUTPUT1(13) <= IN1(5);
	OUTPUT1(14) <= IN1(5);
	OUTPUT1(15) <= IN1(5);

end process;
end behave_SgnExtd10;
-----------------------------------------------------------

library ieee;
use ieee.numeric_bit.all;
use ieee.std_logic_1164.all;

entity memory is
   generic (data_width: integer:= 16; addr_width: integer := 16);
   port(din: in std_logic_vector(data_width-1 downto 0);
        dout: out std_logic_vector(data_width-1 downto 0);
        rbar: in std_logic;
        wbar: in std_logic;
        addrin: in std_logic_vector(addr_width-1 downto 0));
end entity;
architecture behave of memory is
   type MemArray is array(natural range <>) of std_logic_vector(data_width-1 downto 0);
   signal marray: MemArray(0 to ((2**(addr_width-12))-1));
   
   function To_Integer(x: bit_vector) return integer is
      variable xu: unsigned(x'range);
   begin
      for I in x'range loop
         xu(I) := x(I);
      end loop;
      return(To_Integer(xu));
   end To_Integer;

   function to_bit_vector(x: std_logic_vector) return bit_vector is
      variable ret_val: bit_vector(1 to x'length);
      alias lx: std_logic_vector(1 to x'length) is x;
   begin
 	for I in 1 to x'length loop
		if(lx(I) = '1') then
			ret_val(I) := '1';
		else
			ret_val(I) := '0';
		end if;
	end loop;
	return(ret_val);
   end to_bit_vector;
begin

   -- there is only one state..
   process(rbar,wbar, addrin, din)
      variable addr_var: integer range 0 to (2**(addr_width-12))-1;
   begin
      addr_var := To_Integer(to_bit_vector(addrin));
        if(rbar = '0') then
          dout <= marray(addr_var);
        elsif (wbar = '0') then
          marray(addr_var) <= din;
	      end if;        
   end process;

end behave;
-----------------------------------------------------------

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-----------------------------------------------
entity alu is 
	port( X,Y : in std_logic_vector(15 downto 0); 
		  op_code_bits : in std_logic_vector(3 downto 0); 
		  cz_bits : in std_logic_vector(1 downto 0);
		  OUTPUT_ALU : out std_logic_vector(15 downto 0);
		  carry_ALU,zero_ALU : out std_logic);
end entity;

architecture behave of alu is 
	signal OUTPUT_ALU_TEMP : std_logic_vector(15 downto 0);
-----------------------------------------------			
begin 

zero_ALU  <= '1' when OUTPUT_ALU_TEMP = "0000000000000000" else '0';
carry_ALU <= '1' ; --if () else '0';   -- Add condition
OUTPUT_ALU <= OUTPUT_ALU_TEMP;
------------------------------
process(op_code_bits, X, Y)
begin
if (op_code_bits = "0000") then               -- 00-ADD, modify Z and C
OUTPUT_ALU_TEMP<= std_logic_vector(signed(X) + signed(Y));

elsif(op_code_bits = "0010")then           -- 10-NAND, modify Z
OUTPUT_ALU_TEMP<= X nand Y;
end if;
------------------------------
end process;

end behave;

-----------------------------------------------
library ieee;
use ieee.numeric_bit.all;
use ieee.std_logic_1164.all;

-----------------------------------------------
entity top_level is port (
	a1,a2,a3: in std_logic_vector(2 downto 0);   --a3 is the address where data to be written , a2 a1 to read the data
	d3: in std_logic_vector(15 downto 0);        -- d3 is the daata to write 
	wr: in std_logic;                            
	d1, d2: out std_logic_vector(15 downto 0);     
	clk: in std_logic
	);
	--is port (DIN: in std_logic_vector(15 downto 0); clk, en: in std_logic; DOUT: out std_logic_vector(15 downto 0));
end entity;

architecture behave_top of top_level is

component register_file is port (
	a1,a2,a3: in std_logic_vector(2 downto 0);   --a3 is the address where data to be written , a2 a1 to read the data
	d3: in std_logic_vector(15 downto 0);        -- d3 is the daata to write 
	wr: in std_logic;                            
	d1, d2: out std_logic_vector(15 downto 0);     
	clk: in std_logic
	);
	--port (DIN: in std_logic_vector(15 downto 0); clk, en: in std_logic; DOUT: out std_logic_vector(15 downto 0));
	end component;

begin
comp: register_file port map (a1=>a1, a2=>a2, a3=>a3, d1=>d1, d2=>d2, d3=>d3, wr=>wr, clk=>clk);
--comp: dregister port map (DIN=>DIN, clk=>clk, en=>en, DOUT=>DOUT);
end behave_top;
